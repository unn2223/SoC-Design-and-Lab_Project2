//
// Copyright (c) 2023 Sungkyunkwan University
//
// Authors:
// - Jungrae Kim <dale40@skku.edu>
module DMAC_INITIATOR 
(
    input   wire                clk,
    input   wire                rst_n,

    // FIXME: Declare your input/output port here
);

    // FIXME: Write your code here (You may use FSM implementation here)

endmodule